`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5uCSOY/tVZu2gAx3iQ+3cAfre8DzK17YzJEPlnAllmPldMDskKzAxhCs8NgQkQf
HjFF1DLE99rHmp1DfEtv6EiSPjIPU/qe5kd79pYwirssAgAdybu30OwT0wJJiP8X
vMOMKBm3hPVUaLQ+VPsZv1lCbG0FvmdJJsQNHhLCVRgc/dX6xAkxzw1+eQvD7S53
b57hkGNe1ZFu/ZwhqtrkC060nACLsBLV9qi66IQ/4mWrZjidEpiqxPP5l0+55PxZ
afC+S+O70ZmY2zvlF4Mj8wGHkIxuw1Hf28C35u8zmQy6gqKqeE+9MV9MQZUg3UKS
/Lc2Zc3FbRFf8fonJFkt2iQ0sTiwUUp2DfzOTJQxx07/vDVgyYR+JDlAWADz1GeT
1uhl1PYEPEeWYUYzSENS2KrvPNphNm9Ylt4qyDS5nguBFOym7WDQxobwldH1oA5z
UJSqQlVidvrdXzQ34d8aiUYioULFP16vezXO729hH8jDUSIaTxkObxnkEqkKZWLY
wHgFB/x98TMb2I7yoZg/iTU6W7RAEpmg6kR54DSdUjhXxXJDkphjj1PvbcCQm10v
ZV2Z13baS4gHq8mud1PQ+ISqDGFWHFBGN0aLaejCCvkJ7Ub4sdScofy/sw+i7D3J
N1VqMF48lJ+5hl33sonLJ8DePnpNZRPsPO5BBjn86iltrXViVwNl4nXV+QqBFy/p
4oWD4TckWOodlFeNxSHfhIryponygVmAkretZqAtJdUG5LavmtK6FBMdsYo3BKNv
SnRdnGx8QMtIKo27LzMIKw3Ac5dXTPAcHIJGh3uYIb/WZvLsADK9DLlg21r2rtho
gf3ZPb+ABPOawFpNOHMx7bwAc73GtVpu6u0oZ60Tcg3Tbc5vLPYW2IvcHGD1h5t9
rBRWCZximgz4InRVWIQ2/1IKTxUe8a1atw2alOQ2y8GNMzu5L4vY3O4PCwvhzrzl
Rn2ALcxYcjNL6g4i7ZAuk8cDD7ImB+Q8BpotRbP+gnyoIHjC+IYt4Fg77QRj42Mr
eIuREMTshSx40sr4XmsWVVcKGskxxGlJE8OrPpMVg9A4Ko+rD8X2KtNuWRzN2jtx
eOT10yQcgkbbJ8Scnd+Ako5KUreaYDW3SQnyEklDg86JT+SZwZSDZo7Nynzx81EM
0lMuxGZSuFU+BovV6sXEO+PXC2q6fwVMHhsR1o8ncRbLBsvhkIPg05sWkxaR8/4M
fH8kB43hDCZskT4PLcsvqMd04rkdgeIbhjpf2Nl12XiWGIiHaIc8KB70bdgZo3q3
uoEWL5k18DrxiJKR/pt8K8UOxwUYkcnnbVE19YI0RJESqc4ns70cZJzyXyoCCVHK
BPrdZDZjWMUhjuBkYItgR8GAfRvGWxIS79WdLiQL0p+Py8Nmc3SFh/15uFEUHixE
nmDo2xjaVU3sDAuDsIi1Qvjx3NRkOH9v7nCxo2Y6ptyw73r9fzoWJb7Jot35qf+e
Cj4U4hS0Zry7CACN2oowS26izTFYsoYkNi8OcQEYe52u8UHuZqcMu26Tw46XzKJi
64Gpx+d3G3ZqCirWzzQHWF1sgNLN6E/fzi2K36+5kbvS95KRcxaveiF9Ckb8bUbZ
odtbjgDcade9IOGgeq6siAvF97I0P6TNOBdsGjDD2qRSiaPXng72z2IoAFIVMMOo
g4vbwrbppq9A3iGZKlLHrGhzfxwlmlUEhSYOZ9Nr+FVS+76LdpbB2fWeNmrGmRR6
wAWt/IZvhj4SuuIzCQhfNspRIkYRpgmJAM+FitctJkE/HntT2H31kT2LNp8McWkb
6N4Ns7baMdbGchRwPZx9hBp+PP2VaqNQYFTpLCa79zxurzRrRrQwJL9d+CWhdS/w
R+FCxBmn0Nl5PzGiSSEnXiLz3Ex8l0A6nJkT+QQkNrmQdWQkpFvdK5Fr7//Ebc8m
vLQ/pSUY0JxhdtbMP97mnSp2p77yZ7UQTDKZEKAqleyhsX+VeX2pGo62RyjP4WSI
aar6o1Y7zDXucnUL1tovqkU8/GghlZnkV3DtKnGwZJ/W+rBgflPxR7zdc1Y2Cf8D
GSYKBNJVSjnUSIkXCGLC/uaUbsAxIOTk+Fb+zbTi9j9v3kXblXAKJs1zHxdqPtLL
Guj8LDmAsaZ/Dlne6jzTePRRITMShThVnm5A3aKcin+ZVUzzYW7AQXXpq6gPL+/x
lm8LUIqEKtPauulPD4VrDe0o6Jv/xdbwuCODycCVNGEWfYRB6BmO3yb1H70aHDgI
4B07WYdrTQeK5F4Htg1y8lZf+slwDRTb4Mq4mrF4MduW3H5Vcxk1R6w6KnCOj3Ze
8QT4lk3TqRLy+apCG5wHHh5gXgX4yaUhsfdw+zslG/ZnTTCEVETl1cyrqUAaYbr9
Qv4r171sEbeKCG2wAj0dxrEOwpR218StiVV5uFyzc7D47vQtMacey4YSFSnlasni
Zg1sXAk9nbH6M2kfU4P5tOQJDoDVv+WaMocaQC330ltyq7B61TGmc1LEU1QTWPjW
xDL8FHGzGndwUIBISkUeOsr8teLFJ6juhbTYFPRrbn92bvryzV2h9aczOv5C/8ZM
OKSgcB+EeY23R2ZquFUDUcHlTniA6lOMokCZXvsdCIdLRqCMdCZI2erEko9ft3vY
K3YjAgzC8y7IvnpkwF8d3QFBt7FzycYk2v/vri0HtV46GknoGBA2bh2F0Qg+mlM1
W7mjVqh63yI479Ql8q7FbktwHaQiVvuEv80LCeJiwdmnMVe8PG8DL1rjCeFSURuN
xPx287S2pPySCjXoA7prk1D3SrZ3OZqSsKdC7wiVHdcaaml3tG5Jk4vHE9i2MnVo
FsghmsNd7WOW2DQg59vySsByXIIpeZkGgP3noA6kpt4+UwkYdtUDu67oLebzlpj5
Wiq58rTvOjntTypf7spBEQD09iZfoahXf1i04JVomcyor8aa/WhbFKEbfYPLODHi
n4EzbzAJuW8QwjbIF2dufskWopN2tuyoXJueDGkeaqkLEe3hAxTSEl6y5CX96aFU
xatXka4Q51PhuTYsx7BpuhKTB/VgmNYLE023yEDGjXFTLMON7hKgpD6wMTnx9zVS
uiNqmYpq52NsR9VSlmF7Xb0zoZmrS4HQmLjHCF06vDJzWPlhQ0K4rMybpUwpidF/
j+WGl7eHSBC4G9LdwAiqmRbe5c8GAJRbQwHkbvl4GMPlbRxvpxaBbjFBBleMN6jI
BI81ok+y39omsTCXHRJ79ZksshbJQBhgduT7Dm+p+eTghZBDfz62eYb4RD1nAhC1
65idQQQubSMnPz50/G9Df5dSht+RIeEG6wglL496UwYwVShsTzeX2OW5LUgBQk5G
615vzDatkHPnMu8WiEVSXvZxrZmEKgGkXhY4Hnj7EBzp3mXSOWG6G7U3ggB0d9jI
wKa7tsOtBqgNIr6sNhm/O4fdaB23jKz+nPViYitvSgZn6qZqOA8rZhU3yH9fGxd8
GMIyRKTyckDZ9k18cBumCR3MBmT5u0amiyRVzBLCIpUCTGYkMGWt52lhMBkbgf0I
2TFzfyTUtNd/TGanA4uWJ1jpVm12eQ/KWZCS/Xul1KK01KY0zSLCkFFWudfQ40nw
nBECiJ/WkDew3hUhaGzcfBhSbndPOEHgs5hmDvHfO16xhybUBX1O7Usk1Fwy1KN6
RdiFrGkd1JqaUOXlTzV6X2I5V/pxLsZBjNkAIOnA9ylod6ygY2AX4bRcnLHtOtij
ne2b46biX0L0/2UA0Ho65Tdbg61IspeGlBWwYJgljpJhznUxTq+SlF5AKVeCIacD
8X+2OZ8pD8NCdMCGlVgDNqe/0RkvLiKM7K/kJ3mvGFBKlBy/BRKB9QPEifjSSnDk
dQploljhcj9gJp5BMLBGOFsy8143/ehVBLY0M+TM+sTJqDWI/FIMjTv1V/m1p5yg
nC8NskjvnrUihbxTnBUjaQXaGHr9AKIFmVIUzzZuv/tLAaT4foCzbi//5Q1AIjS7
sOa2hBL85LlD69BY35+UtrGhX0pUAJubt9Tq38fGISydyJx0sgnbjfkpAgMsIoxS
cgT8+nLz1qEjV/3/tRom1w==
`protect END_PROTECTED
