// Include Checker