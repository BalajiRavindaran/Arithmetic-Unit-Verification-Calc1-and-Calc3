`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3z3eS5JD029tU7BDheahv1tAizQ4bx6h/lmJL2+TBxb1uemAHMdLWRnXoW8z3EbI
9a1l0yJKTfBPhX8nrfv8bAfvt+3SIUfvzk5O5MSN7uvfFffRA3AoUne2zfM270Qg
h+dYPFLsARK45pYnHIUBSjfxCfShp3N37QIy/22DKgsL2CmuzCGjA/9HDsTyVgJ2
M2q/ZlBW0VqY/GQz0eywuuM29nL8rV2YpxgoFxJr/nPpx5lggKwRByTVikU6YTvw
r4IS3NZdhCts6kGh6v14HTWZb4sWCWhA1srRJLUJbHvIEia1xD3ziN9mDKDdWZPc
LNmHh+SK3VYp538SUloicoHsKo8weKlKW5Fe6uGKqlAbcrpnpmrxzpWSKNGgffh0
TmAJZrEFa1lpTUPZlgsBTjrlmuVUQZ9Sz0q+moX0Kz7pa7njgLjFNZHEEN/XU/P+
sBfGxY8zFFRJHXJTVjQIM6L/LPJeV7WdgseQJPid0HkNjJYqWBwYz/RQfFbk9McH
`protect END_PROTECTED
