`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sqBe7/VNOpDSUuLLxDCWrM1KxMaktS8/c0QijceZCjfkHDPE1ItlXBKTOq39JFvS
cwqD1GYmkLnQkO10o/+jBShyOM7EXo2Pt/dsy6SaTBRVBTz1ek1Nyq7K2Z+/vzEg
vL3SXrMZCoT+0rspAg7l62xzili6nnH/WP+RiartrkPP/LLB9eslRDJA9OvhC7B1
JAOupGcJ0YyW6Z7k9PNFEi7IfuNvRRToGOLamgppPGqbEVQmFih1Q2gCjPSNHhgY
WygowgHE5NWodRoweOGaOLBEmlWMjtVsbCfkwSoxdlzs1bfJtOmxKv3q8QV7srtO
WcTetnCwfUEV2YqktQVT8Fumy9zruveRIkPkagkcL/bgCKKJJ5NUyk2gx1GICBLl
BjKaBGVbPycvpvoOm4xolRZ0VyXmOciXJHmw7Nu81IDYQlILgSWssoWSQm+0iew1
AdXf9NFo5pPf4Fysg3o+vw9PTWKZpaAtbG6yzpy6n3LzRkl4oYIr2rlQvB9GeyK+
ZGzBKA4PS+nWNs+G/I/6ocy5mRQkgP8LIax4ZeSFFgNDiL8Wis6q4ZKQ8t1EMDGH
+/yNmlwXmJ65IrcBOxH0eeWDDsQb3RystimvcYqw8jmoUE6YN36Fued7MOtmf0ns
g078IgtfmKp8XoOMSRU+zVYVmHzxknf/l7RALv2JWcXIvrgLH3iMWOcn+W6znlLn
GkVZj4pi1mh1dIUDDM8fhSckuc7eqe4jJXNStJ1NNUKw3vUvw50ntQvetyp3o3/O
O7NIrmtfEVPIRLIPqClSJ5rNORD590+SURpbhRo2QLoIrtreesndB0gT6cIKzMnA
ekkWyOlK/ZPSPhZHWq8WeRs5kado9q8u6EXjj21QmrAAjE/1WVEuYfJ+T6k4Lpmi
G7o/AApf9CoDF5OFc/lqvUWLjn1EMTIJZOoTznOhlEbhJFfRCsR6svdqKjKzrN1p
VjjqPnLSIBxlJgO1lwFXy1jGGiclymtKNq2kW6bgvH6cTf1HAUDSQQYcoU5wI3/8
EAE0eoP2kh7kI1trkd312wcQ7eSrDVglpKv2It1TgQIbNPtTAH3B2jaznleMDvsv
kXiAWM+Vq7CGy3zzHvzgPOTAfNCD4HjvKWXGio7JHb2UOPUFe7vgrCQrfMLK3pLM
/xqp4yllza3B2F7IG5VPtrf9OqHD//MujrFkVcIpkYSdXqd8smNhBUwf0FweOCr2
ISy7X+dRC4ep+HhPI1xspc12kF9HfZjK6hT9MJXSYYgzk5VzzLmcrlF6tG2sCCJj
XFGj+WAUK5PzOCfKXyiVBWpHJfHCTu05aNsQUqsGr4+EA1zJq9+py0kwwcyarWio
ZtzWOE0pA2S3yt0DMsEwsTzuhJ/y1nvBVGsaVKXtHEHRWRAuJR4PnWBY88N1EZpb
sIogzKYk3LhHICSkxWHVdrOKMQJqlkj9b7aVh9e8gGRiHxM5XkNjKBXBg/h+xJay
wY3HhexPF6tZ3vD3Y65iFyulfVG9Y3mi31K9uew3gfZUnFpbrT5gIafNymU9l9QE
ZpDhUDfA/JTZGvljx/P0UGt3zQG0ww5GUdCu/PNWtDj8MpS2pTyvFBui6rKe0NwJ
B1yPjHXah3XXBzMxeiWf3pZ9eLWwXL8jX9nmXCl570p70MlPztw47KRv9F1rvshv
pmV9CzG9qUwS1t9TTDYtQ6baJi6Zpu3uge5j3oo1knBx1/SgderomwHR43ubuP5P
OskozOYQijkd9NAampO8ZOVo6c0ijVKO2FlCGFM7qS02xhZ7vuFIuBFUOSbC8ysJ
DmTDb1TVnRrLGfkK9bTmU3+DQlc00fet1AAhmSy0hQ3UtOhEvL23VrsJcgMkobAM
3/630XQDrnRZznjl5T1B/lGTjrSzp4N/Ypj+0KdnjCZ0oT5mMMPUV+ZtyIoPUTpc
BMlVmCFF/22Q/TlsshSPGTzahxjYPXyY9jwxzpGXgMBDmeGDSw0dZvVBU+duTAyO
l2drkkttnsGCuZsWAFQYoVDux/jplCYu6gtGHjUCOWeQRv/sYHZXYJSg+oX0D02i
wNnrPE83nLalYyq549xuRNfQN4RnmtY2Rhia/1WhWWLDuMn7NOvY0r6IcWkqPZPD
kpFVW+gkJjz0oCAcLkNyj+Dbjz0u8CzbEHns52G1PnJJA1UYvYzBJfugmnOJJg0V
1IR0bbCketMgZIQin/9BjCEKxURM6J/SXV/QmFLre9w=
`protect END_PROTECTED
