`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6wSlYg65iOZ6vraXUUKcddPqir3UQO++cyin3O4dcDUYDu7u9q+Tjcu5U+ZybqPq
2h+VZfd9Bp4+kLD8OUdNVaOMjcgPZTFQ7ESDGcjInVbuBKA+J9jmNoowHOyYVi3O
dBYNoL1EjJ0Tuyq/OJzV+BFkdlRjTo2h7tHU50Rw8nqYZ3uRV68j3NL4ObvKfMSh
ELBGbPAb82nw4I5gaUmCPTuHVBAJV1ztACX9L6JANiBhvkYoDyn6Qcw3pbeiiu7j
lURcv5WAgrX1QGEVtjLu+rP/fwYwp4OGDG7DN7qhwoAblol61HkoJP3BMzvn2R8q
A3xXtpt0r9nISdawAUmz/ChyPq2ehp7DzIJE5kA86yvmZnuOsWGscZt/jE9Q2uPP
SnKnAjPcO5yimeJ9qb4kNN0DYD0oHXLJXvY2Qy/Y4j7nF5rm3mVrXWdhKnd/HhYu
I+Y/xVkvYuhBsjnx0jcdizslM0AbVXUf835OAM09H0ukO8yUUONzc1e85S/F2gck
eB0V3ZLIJXioWHPzI9Ed3/D02hmkhfp/vd3UIYpghyAwKvOdYBxNMxDxqER8NeWv
39BX8A3EhzpiOu1foXPOwHO5nUH/KUTZNC0dTQYlR2+IlenDT41fsdHWI02w/vlx
FmEnuejrK1gn4l3pDCP1Yn86uW7Wn09Q0IWIPXe9AonCKhFaBQYH7YTXhrqtkK5K
S0aaGQNOTlJZDMYeb42AONKYkrSiLmgEDSid4X9zAakzVPyTOrqCHjGV23Iouvy3
rfwcwr5kslxvevlJT7blVoxYCFlYzbTFcd3u5sv/abUvjszJDOj2wC1mafPoJ2zy
n8+ecHGf8vuVlItUDO+WObGp6Wh80HvUFpaCGIbeir9RTE9jHzQ1Jhon4Fz8H6lc
6jBC6ddSNjNni8ssZF+h/DPgzXWWo7XQYbXL3uklSajoIZMlHbdHJ6+PTQ7orKhl
fklr9pjc7jSvtNw1SP3SInVB/qpSaiVSt/9EHxQw91XgAQQxvOt5/gBGBFBMz6y5
Uwpam+pCUGRRuEhLtHxJoyz3+99aOGH1ljBYMWeYB0IUtuXxjHYUR5B/RJcc0+aM
AB/7nvYzEO9zqO5U1J95S2TkFySAUC3qBV7326EhJ++20AR9sI1dA8npHMFgRaBT
WXiS0SukRp9dohVZijtiPALc2u4WmuOTYBtOpYDcOmH82aqmmiMLRPIw2ix+LJPx
NawrkqLi4iDRIZTNQ7cVVqyCdOb2n9xmdQQDZuddxUictM9zu82CjN74EK180GWf
L+ZVz4ESjKqXH7dhjw4K8l741etJxOf2V8hTBzVjGByg/zivKskZVO39WJ0ZAd1P
3zgx+zQNnOZM3ofp37paJjkLx6F7nrB9jvBmELyWoPYSydEHbC1/EG8ji54U6LIS
8kydhdRrmyFjJ9rI+WksgbZ3UeTViOMk++mmycUyyZ30shW1HefZZk6eNYjubrMg
ldvCKez6IdWULHlCLO6xTgTnI/3ROxGAC/8hPgqp6gDB4K3ixtoOOq4wqSKJ09TK
V7A2QREKzWGdJKKkT1JrlN52gFybiNUWmWDUG81so32WuaeuI6ormWnFjX9wod7y
u/A8ha0T1wiGj0V7Jj6HOz7xm+0YQPA4EVs8GxozuF6T1t2I8TeNtjNMGgLx+Fur
5mdEaWLleSu0792eSeC/z3HYXIuT18X3DoDh2rUOV3icjVw6/Qki4YQKUmHmYGow
`protect END_PROTECTED
