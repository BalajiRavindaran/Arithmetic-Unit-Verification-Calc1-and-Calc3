`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/OP4SEqlu7Rc1jjVdYc1qjktObg254gjq1VX9FVlR1huKfvDjUM5G4Wq4/BoZVH
zu90wWZ46yYE4AXj8hErfdM05JEEnks5rGqrZ5O6YY7tLXkDdtycv8vbvC3NOaDm
95hRFurtFQKeHuVrvfPAIaA1NjAIq3pmMhpMXEvES5tB1bnAfSyqOYk+cM4a2zNg
BbhMwby0VueMbdYoXzjmXxQXDS05nSHJEpM+w9imvoicGiB5gnEu+egaPjvq0BWR
LdD0G2DTh0flAcwCLGiQEv5H6GVkxJ5Ln2u9WE+ghO7iLymqtBwCWHX/qM50bM9L
wY7rhu7ci9ZRJLg6m6QEQhmyAmV2P9X5JWzH9x+KG27h6RN+gavwRKNXopI9YGJK
j/36GrxYfxZ/35fiiWOApED6ydy7pWXkEsHwlTWyj7fWKhpHf6skUmwp2VFedVXa
peo+9HKANH7GbokTYx49B/uMK57zRBcDxRC/27zE6Om2/CeOQyE2fbnOysy3iDsw
Q3MmTEc4NVBryupR1i21g3XkaY9EWZjuS7G8tcBQDQVGw+FtyCMMruVETk947mJN
VM0rnbvFgdI2c3pUyVEhWtix0oQ9ffRysRdF3Vra8VKO/jz0LgAfsw/jtKFgkYmm
sV9LDhfGPyOgcjvDOcRU/zUoOUAfeLeWudKRN27XftRBraGRagkZ0zdDEYGZRjn+
qPJA8KFSRa3GZoecIeU8ccCKGPe11UHs9z4vh22nm0yRjgQ0edWY04oUFS1O3AaB
i9SsH/SSZnL6ENgMyByGkLnAiJkkrTpqev9HneW4ZVUytFA/xyU4mK3BCCTII88E
KImJV15mvyKBC9KbcPKRGRdY/jKnZvdn44MLN8uHfCS6IW2hwvZQY8yyOO6h5I/2
VTPuihQiUbznPoSIqQpAKY87tgl84ROTEXEvfBvG+cjTyhqBqbZPL1jigz2mhpIn
bckSaI1aljuOLGbOwMNcSVBtr4XhV+D+kgBIj6cUa1OgvtKCes0CS674gmy6XeNR
NnYzaNJ5lS8ssFgWyjyJjsM3AicroUAei1RCD5IpbQ2EKF1c0OZOteJrJvKA0R+d
brD7w+yyozFg/hekMA+gUWHsY3YUqZ8agXTAJXhq1qJMnn10/kB8zPOKgSWSurI7
CCLcQ2yJJKlDqOtFI7JLwItoE15PXDCY/7lfuwXO/lgu85LDlgDOvdiICuq4u0UY
CjfFp3fsvgaayt7zuiTQjb1ciZckW5hu9ETqvkHG3G4hXgUAmBfGIHm9XDi6IHCX
s0KrGYKks/TIOTaSncdKWYnE6T9aPmQRRex9L7wJMk5FujDIdsUl33HL6KOMcsyc
LSR8BlgctOz1O0iXacsMG5lRTR+xmyxR3BGFPxJSIPs0YDDWOzsZGTdhx2mtR1s8
2dfe7Wh0B0dvbDX0CZiVVJJrqpzDkIYJyWBbJ1OBjOBEXX8rScqk5dEXF6Lf5cZA
lyVSG5sqyuz1BLFI60PrGyBWWVlRq+/nUp1aLStq3XHA7CywnGy8SSUR+H3a10kl
6n6hgfux04aZyG0zSdGWZMMQf/R2wvYIjo2iYlbgpSQbe4lgF8fb4ceuDMQKW+ca
1zl7hja81XW57F+2OOpVCb/ilIjJ5hJm3qs2u/7d+BM8OulYCb5TaDJswBf4ig4l
FcG6w3Oy0a9zyxM3fzZ+kLFn0FetOgE6zUElSpCVJpjwBeesYaoLRAujrRvM3n6r
dKOKnhCRxX7T+eKk1KVG4mBitJjEPJLCGdq8zTw+toysCAVcd0golfSD2YaZhR0U
7vjLs/Hsc1oZk2cDRdYOjZH6TWvhZahHoMdnFqw30zrMKasYt0kGZroehNraCqLb
5iLvI3BazxO7GelrbWuzGZiTQJqxbgYvrdDzcfxxD621QH5DdMZKqObM6wF4ecOQ
J8nqZH4174ICX/VeMIiVuQ==
`protect END_PROTECTED
