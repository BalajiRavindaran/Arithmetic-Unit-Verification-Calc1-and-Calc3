library verilog;
use verilog.vl_types.all;
entity Calculator_DUT_tb is
end Calculator_DUT_tb;
