library verilog;
use verilog.vl_types.all;
entity dut_wrapper is
end dut_wrapper;
