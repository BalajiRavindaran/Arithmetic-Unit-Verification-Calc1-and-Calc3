library verilog;
use verilog.vl_types.all;
entity dut_interface is
end dut_interface;
