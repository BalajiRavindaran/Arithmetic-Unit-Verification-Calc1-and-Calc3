`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
355EujoSM6ZFMb4IPxdGcw1Mz+pVDDx3Y7siE5SkopMJN3zaJE3fevIbu3rP611f
tX+/68iP4KShDZD19fAVun6OJW0InB/1k/ol4hHmcljX+ar3QYH5nQVEcF8Og2N4
RvYyUfK3uStmSdbqjKtRhB+aBJia/Mf5ao0Sxq199LZcEBbdCrB9GpsalEoLUusC
8zBGYgwk26nyNMaXWUUbIVEZyJSDVvLSE1be6buC7PDLZf5AEIsGoYqQViMmL5+Q
PZdZ++cxHakWX/kxFFvGZP945Hod3CtNRtQ/MKIAOXv2FmYLQ2eNSWKjcCuvFZiU
1gqc7J704cG6ZdlpZfQm6EeJ376+vjjvRJMayXOnRNmB03ZsksqG+TiwbZzsUmoK
ihZ8vH9T5W9hm87uRFeKQj+fVWZd5ckUINREbX1UOO+/dJtNTTXUQcVGazA+xo55
dMNHChQhehsd6FFrJFwwabOmeXsy1npniAwuIMDVECCVXOjZdaTAZvde0icvpAzo
QvkW6zlxWKZ1T964ty/4s+SznkjDaUUy690pdMr+iCfZibDZtIkPkXl0LoToYU9h
3WgFvKT7y9a6fsp82k3Kgkfetgp08Tojd7OtBkyURAVT8L/mCMfE5xCNe3G6Lefa
vA98La90QKRU9EE9OY1aEUk2IEvDHs7hddbGg5OXzlU8cHgGlmoc/U0GSqz3NPMb
SlnPMl9DlAyjlV2puuPdBLdKhJygHG5vQBEl4V1TqyZKOx6HppcXBDIbvUq2I+df
nRGrOA/1HTvuM/L86sy0n1/l6C7hp1oKxxw5+rSg92tsW2uua4uczHAheGuWsyUD
zlkjJ0VeS/t1Xg9z4wkt9f9TxWzUcGu/G3KdRuARfPvAs7n3L5giM7c2x0sv/vCc
fsMjGH1DjQHllwpPkU3a92inMFgc8nT/IFZwdiU6ZIS8Z4IGOfGDAsY2EaR2V+hj
tMboFm4rckdRs+2au3h/rcQuz83/nw9Js2qIbrOTkNNubDyhj8fTqyUblA1Z4kgG
F++kE8W068GqeSI5fgOV8NRJakTssEEeJC8fhe+MV7460gN1KE2syEykKk6/794E
5aLO0XqeMm1pNFlkIuJKvvJi6H4MyKfvpiIgZoh2qyIGaTYw5QEny8z/i/55KNyY
AfumugPeP1xLnUoHMSScYYfybLsVGz4M67fBiSAA6QjM0HqfaigFi4/Evz+iUtG6
X1e9C6acnB5rcqPUlaToQsgRHvolsqFKA8ibgp1YqElyUXI+FEY9NGZfVAVSINEI
YgQv6PhP0MjYESUjkbdLZvH0PHpkL5U228NDxcBYAPhyzqQitQK35DPnvdp9o4gS
sOb0CvRHEJtyiE8kdMkQ0MGd87w+ht2jNAYIljK/bhLYl4tZm4IMvOyPDJpOZD1Q
cOLr1PWE5k4gTfJm9X7/qA==
`protect END_PROTECTED
