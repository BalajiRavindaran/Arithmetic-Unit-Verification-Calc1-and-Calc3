`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/iebAAPT0VVZvzms+nWsxlg/GpHC82XWFwbGXvMsAz6vM0JboGYNnvrhj1wH4WV
DTqxBg9xm7vDjoQc2YMmID4psRcsUrxq5iqFpR9D8h0ZH6X9m1JdbtktO1dpbv9a
HXMjh6BvgOZx3I+ZNUrA5sOKFIbB8b09xykCCdlOZaX/aVp4rbbhkbad77+3f+gF
scVnEuMOmhqlivUYmLmOsO+8dKmw7Hd1o5ha3wN7Hp0HoquyoCLrNdVH28hTZDch
/4bw4uhvJgoyiHKfLUm9AONFGuBvm3oCIBL7kVd8YYG5yapK+fklJP9PRiBWVu1n
q7T0SZl0MYXS6wUc0jJzfl/l7QXmAFnv6HpyAwxLC+T2j59USXJ6nKJprATjmphM
680NKuUoVOCrz7xl3uWl1fyQym3xnGjHwhUMZEpgQeFKb/W5RQjAxQnxrpIIy+JF
Ui7g2Y/vmPrqJ5uPDyxqpFksrYZFDLQjqJ0oKTastmdy3oHZM5rIWKRctDtzzzop
xEwRfJlckXmJIS+BB/Rp3C/rfTnNnmd5mQM6WyZVMxWRORRj6pJT4g/gQUjSQluR
foiGasuAMzDybL1hqTRJ9iPuRCZasHJWQWMGqnUPQGp3IAFpnnRWMCSIC9osZAaC
NHOnoW+sNubohXNTeI9f4pYJno93nT98aJfAgEym/TWHF2vPxpYtc6xwn8peUc0z
8GEbx7VWc+dy3Bcz9QETuSaLde+Ae7j6IV4JBsBWE4y7f906g7FU05cYbOeQ6Z+Z
UFvDAixyKh+9/fpnJw2DpmIuOtsiqIRS3b+LkvwSOOTpnfJNwQaqGhqRV0hvF3j3
+gjJqtL+p7vAzSHoUat8Ken55lNukmeiQkiDt95h3tOZ9gRiUmrZRqFIZoquYY17
Q9LOk8SNl7rWLaLGaK3gYrWlHwzkcMPbkDHvDa5QvWaX1MmRtif7nff5qCZo4z0H
ShDJc54m0p9nLx5P1D67CMP18gLlA+3AO3WQ7V39A07CP+DCMyxEb/LWH0s2FsZ1
IyOOW0J3hlt69FCesg2AvAg/cl/cilG7Dh5uNO5CymuGmbIv+PXHyPeatTmw6rpB
HwtUogysK0FLMWJs8JICMV8vvS3Gi1u/Zpwk1iFuNvvXe9B2fksrBfwojvc+WFqt
hu6ruYVRD1kT0jjsPkSlDrtzRp8Q6Zar8yCqXq0ocArmhh2MSOULbERM0nCa1LN4
tx/3IIyVKIy4BMwJ1umohFZoHmr0QQzupN/qvswr7WL0D0Ahdb7LLUP3oYoLEd4f
E1wPoRuPyhaJxnNQNFkH71r+/A2Fxt2W7S+8gJv8zIbD39aS+CUeorIo4h7UyfQh
/vw/I6Htl1mN3/PcsyVXtyEK8SJWEar6EF0kor/G3yCJWwLgRG9iIloxu/sqhsMA
DVFkPk/a9k/nd5ZKLKyXgIHCHweQ8scdBFq40GPqsPM554kzlt8aDkDnDO0US7xY
wYHR/ZPJbdXw0uKOPHYBRMaxPJ9TEEOyb7HL78MLJxxNZ7uMFhU2Q3owtkt0NYdV
fcbQmU+thu1f8SW0AoxAOmV1WsI9Z5cU4JRZrv2+O5UMdf7P/6EXhCmqG9iEZ5/8
jjmTuN13GNE7wxpLbEbNhiPjmwjfJIpFlBzeRlFTjIBvwPs3MCWxlYmlu+nxgLyp
ZecscnYgduAIF91n94cHfQ==
`protect END_PROTECTED
