`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/OaXkBp106s/RT4xuseQCzUYvhDijKEEriDD3MZrhcYy/9JA8SB2eJBq11KJD21
bzEiNzeijpujU2mOLRlKnuXzxiM8nUvL7QNIandX3O7NYSWcDhLpf8ijsfk+j7jJ
+Tkxn0hKYCEifh896lvxFNGqaco/ex2Obi1q6SUdRWsN5UUjXJZTxKa+/MNu4cQC
C50p9OpJfMAO2ZMrNkRpFy7+PmOPYuNqP0X4dvYwkej1v3LK8Qfi2wlDpa0cM3dp
wu3ZbSwUxLG9OmjYR8XoJzdPc6Sy5/hBQjUQmXudFKvvUwgBCw9RmnYefv67W4La
croBA+zUdp98ZD7gmo+p18wsTRl1r5w7KaaqP9delAv+4KWubDtsWnmep66Fe+DZ
Xw3SRlaRdwDrIXsaPr33sLg36IOnN15qaEfj+zPP9DsloO+V9E7Xr2iQjV88U0cy
rZiNQ6O+E/Tr6XO0T8PGj/eRBzY0lrHmqw4rVuM0H2ZMEMBfywlnNsE+ahPY1/bF
nRVSmEzXEshFqzAzK2QQkTaJYY44VHPCn6M96nhI8Q6fxqfu+9CwoLsVMYK6tnir
9LsTmDQZ5TUJth2GNn9fpg==
`protect END_PROTECTED
