library verilog;
use verilog.vl_types.all;
entity Transactions_sv_unit is
end Transactions_sv_unit;
