library verilog;
use verilog.vl_types.all;
entity calc3_dummy_sv_unit is
end calc3_dummy_sv_unit;
