`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r79HF1PnYq7dnrhvRk7hPBIL1E4NMBu58DlcluHNMcvwjF8dqR1C84XLC6H8h57B
aayRcwnhuITw1Oj/2d69elp1Lw408VnJuhyYKtwoEQjVy/GhliVqlf8/m1SnanLH
XZKAsG58xXcw3wl7hk6DDTiw6n6KIVcXncQpjc00WylHviyMvGDqq8XAzxzrX2Ab
GDdGLrhyODSldMVdq9IOoxtDZrBr6dRhwfllokuI+mBtFW65eSEw+woOGsvrb0dL
6SrZwDXID0ec0D6iy3yt/e4/c4LJ1HSeEx1O8rmcbzbMvnlDR250ngPbR+cS/9uB
oAZniQutMVgYjdK9ARkRWEhVQCV21F/66XCi4EdxT7y6kqZaTxk77kjE7QO5D0R6
Uae8XdKALJkmVML0w+fOHXbIvfBh6szVvWVd14C6dtyNM+OL/BHmUD15KO+c7euN
c6V+x1fkJTtDr8Vk1GQYVPRCE5wInmVnSJXsK8kymwU0YVOgSAqKi/54R1EhB/gY
kI0pOpmr4UV2AwnVPSlxuK+HbtS1n1/xS9xXQq1qBmqGHb8xl6iNl0MoMM0WKJM0
UQyk7ZzxAvma0/IcB485sd1mKaLMBi/mapomTRzb9b1p+fEP5d3hN/16Pj1+/gRm
RGCw4hflo9nkF1rKSjN3SZGu6kgvmLztle5dq830BO8kgM2LUxMet3EURk/rz2u4
lynyEanlfch60Wnlbu/tmDytllxAsuX5QKqKDFuNtaJczzGWctfV5+s2arRQ6VxU
Ao4qmrzGLPYlqj5lzywQm2lSjY1AucKQjaXwSQMoT3bWeILY8sJGJY4HzEJfdgwK
zgL883aeQKX0mqu5Kl2kndMDyudRJOaKVUp3WJrzJy3gFOVOKf9VDvu1MyIMVUc/
Cv5hxzpdZmhWKKzgAs8q3ibfD+v5C9BzXd8s7HXg4Z72kiAobN8CTTWJITPcYqm2
DPV47T3DNR0bo0TyTpV3ayyqzbWt4813Zix0gNfPZpf6CJWTMCtBaHUwRms+YUbn
IMN5JPhAWC1muXzsGizBj03etebSZfULaCEicH6OagK0ieaE17z52jWJwZ/2iDVa
SOSAJ7LI3DsekXI4LIvfaCNAVUuK/7HkoiR1xtRRtCBfNN/OLu0UAj7qjjD2TOn8
WvKOdkwj5HzunQCz+tLoVSVoq7wjEhUvuK2z8EaS0Mof4wBr7GS5UksbFSeK+qys
l+TC7zqySmbBTTSuo65H00kKA3E84qz+LrcMiwt0uEtFuuveyDKDbyTkSlpcE6RQ
tCYSGAGhdGb+WWxSdBcQ1BX6z1OiIzx1DbnhUZGTx/E=
`protect END_PROTECTED
