library verilog;
use verilog.vl_types.all;
entity TransactionContainer_sv_unit is
end TransactionContainer_sv_unit;
