// Create Checker