`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mTFuJqmhLFVpbT1vyJ5VaXCM9gSHikXdCXWlaQmjG8/7TosTtQ0wbHIYYMWNIFk
GolgmEb8bx0g3s8zmwvooC4N9SVGKdImxhvvhs1tZr3QdyCVWNY/K5FicE1Q9FFJ
OOUUnla+/ntMq4VGtF0krCAHZ3CFNgtO1J/clJrFCaWpdyT3PeJYB8/9wdDdziHW
+bd3471iW34KuFmV3y6HgNXHbQrJwFpoYY7NPF7giDl55xRf5dEnEKU9wyKzZBuX
RWORIjUR569pLsBqim9uom1qlewceNU7Vte56U/Pu6VORragkuSe6xu79QBYTQqI
H1pkqOIMnLf6lMbuKurp7BYQX83Os4cg7Jv2ppdua+M2ty2rIezOV3a6P8seywlQ
3mm9FSqrIoRorxeNuvO1Rfc8ZvnQmJt49mDyc6kS2egprk3W6r3L5lv5VuD2wgSX
7mmqhMev2trg6QF6t8vrrbQaT/DlMoQrAjDX8rYtkJ/qP+hr8gUDzZmd09+z+xcY
7+tmrSGP6dSAMCx0xrRTgvMRTd2bY/PaQDCRc8nS6dZbCsS8qXDJlJsdoWX1+FkE
y5uFKVmv5As+tfZUcEeV/lYSNb2lRSRgjLMBJ7QWqfP/JaIbFnlifubNOjHbMjCi
Vy+JLeDZUZkIsKuphRZRUdepouAwWRTh6h97tGDs+8E7aS4HBekV5mfJVAT07Lcn
+7urVf2evLrTmx0QNgqD+I3fJXqP3emUXaalIuikxfjl0eZHyb26cor24sZY5QcE
lf7WAhtaQg6RL2XrYTwJOCxfHI4Teh7yc5cCnLgOJCf1gDnaKuwSm8PPGDPwd1bO
/nAp7/IXAoSK8Kz9ltRDvJw26AOgnUOg4NMCy+u3AvIwhxbeUwo0t/PkLDU0dJ93
H2egFCi2oM3e8U22YnsdnFIRC1xhrvsVHhZnP5kUmeWJ9KhQGrFiPEA1clDBSbH/
U16c1zCe1wMQ84sWuWKjmPZVf0/5YEEQA6lCxPIpaqiUAQB6hYmuRe25TLFMVSLa
QfEnFHvZT368AE0M1+tSCb5sxyYdMl02BLT1UuTNs0Li56mnyHokpTcZOlef4Qwy
Qm/nf9PhyaTC7u2Tv4Fo7vtxRJF2AEHNhSGEdeMMsmJ6RgFTDiFvFE9FjFSLdA5L
gAGr+5T67GM21kohyg+chGqCF6AiXPvY0JKUcwr8EQiGpiDS/OMwVbEJrleXRilR
Ga/emYHtnF6uBCrji4Q4u3i85TgGOLL6kAiAYZVYlzzAXnyhqJRky04wyRvkciuu
Aqzgkt+o3T1MVGtgmKs81rawIFwyUMcUjr1PdQX9gkKd33ZxV1sYdyFeDGukmFl0
ytrrwLPy1g4uuSoL41ig3HvSza//Byp28gcK/KSJ5IW5P/aOS5TqjvPaHgBdud3c
0LVLPTMkjkR+TlJOweGYWDfdx7iaUM7ZxjdnuQffKzN5tN3WM7fwPR5IN46vX1JG
2+N7UCmnhzMSgcMiodAehBu7WvMgLS0zX1k+Kp9e5iQLhcouUAKrd6EAqL2X1d0p
c8amwJwZpasvyBQyhE/4WtUpMgzfTudT5HsUKq42kHIyiUyx+F6s/RdfvJM6n6vs
7deYcQToAUoDUPM8DR/KHGf1iE+mJqhmr4i3HL6wkpCBI56xtCxlhyDspLiRc8bv
35CIFPG7uGHpd31LW7q1yNF+YhjIoMeIST1NlptaB9ERH4M+q+Tk5l2ZgLWIOljD
wA0mIVKfBRbsA9vPrwYvWkLSHanY9SG/3uWSHTdoKm3mRmmkiLfWwlLeEpbtXV+g
IpkyRQlEl4JbNUW6YYcNCTpa1T78MWdquTIw+EfOX6pydO9lvl/MPW3BhSegORlL
e6acOfMiSh0TU4GxR29x+yBUfamFfXm+WoLK2jaUjdYhJFtDxiVHcgoCj1dMEHHB
mH3PFdAHXJwEa71Dg/1JDTGi0QTgisib4ljIpVbeMyboBPCBS6NUkF1D3c75NvIC
EokFBVKmHbcGQG+aNGPaTXo6Y8wEaermM+oDdGdwXHrrsO7diHJBzj8PAKlgEWax
jjJLZb0X9XiZJbm271OSpFcaavbY4zVL7S4c6Ianag1GgKti5KZa3nxrBwTjvmQB
46YqsYxHaUVwR/AvqYoh5kfari66YxgSMKTrabyWvx0=
`protect END_PROTECTED
