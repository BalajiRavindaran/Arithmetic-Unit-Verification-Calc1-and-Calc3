library verilog;
use verilog.vl_types.all;
entity sequencer_sv_unit is
end sequencer_sv_unit;
