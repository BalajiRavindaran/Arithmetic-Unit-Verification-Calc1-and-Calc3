// Create Coverage